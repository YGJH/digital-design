library verilog;
use verilog.vl_types.all;
entity tb_final_exam is
end tb_final_exam;
