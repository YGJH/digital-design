module SevenDecoder(
    input [3:0]A,
    output [7:0]seg
);

logic X[6:0];
// 0 2 3 5 6 7 8 9 10 12 14 15
assign X[0] = 
  (~A[0] & ~A[1] & ~A[2] & ~A[3]) // 0
| (~A[0] & A[1] & ~A[2] & ~A[3]) // 2
| (A[0] & A[1] & ~A[2] & ~A[3]) // 3
| (A[0] & ~A[1] & A[2] & ~A[3])  // 5
| (~A[0] & A[1] & A[2] & ~A[3])  // 6
| (A[0] & A[1] & A[2] & ~A[3])  // 7
| (~A[0] & ~A[1] & ~A[2] & A[3])  // 8
| (A[0] & ~A[1] & ~A[2] & A[3]) // 9
| (~A[0] & A[1] & ~A[2] & A[3]) // 10
| (~A[0] & ~A[1] & A[2] & A[3]) // 12
| (~A[0] & A[1] & A[2] & A[3]) // 14
| (A[0] & A[1] & A[2] & A[3]); // 15

// 0 1 2 3 4 7 8 9 10 13
assign X[1] = 
  (~A[0] & ~A[1] & ~A[2] & ~A[3]) // 0
| (A[0] & ~A[1] & ~A[2] & ~A[3]) // 1
| (~A[0] & A[1] & ~A[2] & ~A[3]) // 2
| (A[0] & A[1] & ~A[2] & ~A[3]) // 3
| (~A[0] & ~A[1] & A[2] & ~A[3]) // 4
| (A[0] & A[1] & A[2] & ~A[3]) // 7
| (~A[0] & ~A[1] & ~A[2] & A[3]) // 8
| (A[0] & ~A[1] & ~A[2] & A[3]) // 9
| (~A[0] & A[1] & ~A[2] & A[3]) // 10
| (A[0] & ~A[1] & A[2] & A[3]); // 13


//0 1 3 4 5 6 7 8 9 10 11 13
assign X[2] = 
  (~A[0] & ~A[1] & ~A[2] & ~A[3]) // 0
| (A[0] & ~A[1] & ~A[2] & ~A[3]) // 1
| (A[0] & A[1] & ~A[2] & ~A[3]) // 3
| (~A[0] & ~A[1] & A[2] & ~A[3]) // 4
| (A[0] & ~A[1] & A[2] & ~A[3]) // 5
| (~A[0] & A[1] & A[2] & ~A[3]) // 6
| (A[0] & A[1] & A[2] & ~A[3]) // 7
| (~A[0] & ~A[1] & ~A[2] & A[3]) // 8
| (A[0] & ~A[1] & ~A[2] & A[3]) // 9
| (~A[0] & A[1] & ~A[2] & A[3]) // 10
| (A[0] & A[1] & ~A[2] & A[3]) // 11
| (A[0] & ~A[1] & A[2] & A[3]) ; // 13

// 0 2 3 5 6 8 9 11 12 13 14
assign X[3] = 
  (~A[0] & ~A[1] & ~A[2] & ~A[3]) // 0
| (~A[0] & A[1] & ~A[2] & ~A[3]) // 2
| (A[0] & A[1] & ~A[2] & ~A[3]) // 3
| (A[0] & ~A[1] & A[2] & ~A[3]) // 5
| (~A[0] & A[1] & A[2] & ~A[3]) // 6
| (~A[0] & ~A[1] & ~A[2] & A[3]) // 8
| (A[0] & ~A[1] & ~A[2] & A[3]) // 9
| (A[0] & A[1] & ~A[2] & A[3]) // 11
| (~A[0] & ~A[1] & A[2] & A[3]) // 12
| (A[0] & ~A[1] & A[2] & A[3]) // 13
| (~A[0] & A[1] & A[2] & A[3]) ; // 14

//0 2 6 8 10 11 12 13 14 15
assign X[4] = 
  (~A[0] & ~A[1] & ~A[2] & ~A[3]) // 0
| (~A[0] & A[1] & ~A[2] & ~A[3]) // 2
| (~A[0] & A[1] & A[2] & ~A[3]) // 6
| (~A[0] & ~A[1] & ~A[2] & A[3]) // 8
| (~A[0] & A[1] & ~A[2] & A[3]) // 10
| (A[0] & A[1] & ~A[2] & A[3]) // 11
| (~A[0] & ~A[1] & A[2] & A[3]) // 12
| (A[0] & ~A[1] & A[2] & A[3]) // 13
| (~A[0] & A[1] & A[2] & A[3]) // 14
| (A[0] & A[1] & A[2] & A[3]) ;// 15


// 0 4 5 6 8 9 10 11 12 14 15
assign X[5] = 
  (~A[0] & ~A[1] & ~A[2] & ~A[3]) // 0
| (~A[0] & ~A[1] & A[2] & ~A[3]) // 4
| (A[0] & ~A[1] & A[2] & ~A[3]) // 5
| (~A[0] & A[1] & A[2] & ~A[3]) // 6
| (~A[0] & ~A[1] & ~A[2] & A[3]) // 8
| (A[0] & ~A[1] & ~A[2] & A[3]) // 9
| (~A[0] & A[1] & ~A[2] & A[3]) // 10
| (A[0] & A[1] & ~A[2] & A[3]) // 11
| (~A[0] & ~A[1] & A[2] & A[3]) // 12
| (~A[0] & A[1] & A[2] & A[3]) // 14
| (A[0] & A[1] & A[2] & A[3]); // 15

// 2 3 4 5 6 8 9 10 11 13 14 15
assign X[6] =  
  (~A[0] & A[1] & ~A[2] & ~A[3]) // 2
| (A[0] & A[1] & ~A[2] & ~A[3]) // 3
| (~A[0] & ~A[1] & A[2] & ~A[3]) // 4
| (A[0] & ~A[1] & A[2] & ~A[3]) // 5
| (~A[0] & A[1] & A[2] & ~A[3]) // 6
| (~A[0] & ~A[1] & ~A[2] & A[3]) // 8
| (A[0] & ~A[1] & ~A[2] & A[3]) // 9
| (~A[0] & A[1] & ~A[2] & A[3]) // 10
| (A[0] & A[1] & ~A[2] & A[3]) // 11
| (A[0] & ~A[1] & A[2] & A[3]) // 13
| (~A[0] & A[1] & A[2] & A[3]) // 14
| (A[0] & A[1] & A[2] & A[3]); // 15

assign seg[0] = ~X[0];
assign seg[1] = ~X[1];
assign seg[2] = ~X[2];
assign seg[3] = ~X[3];
assign seg[4] = ~X[4];
assign seg[5] = ~X[5];
assign seg[6] = ~X[6];

endmodule
