library verilog;
use verilog.vl_types.all;
entity tb_birth is
end tb_birth;
