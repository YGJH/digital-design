module test(
    input 
);