library verilog;
use verilog.vl_types.all;
entity tb_fourAdder is
end tb_fourAdder;
