module RGY_combination(
    input [3:0] q,
    output logic [1:0] r, g, y
);

assign r[0] = 
(~q[0] & ~q[1] & ~q[2] & ~q[3]) || 
(q[0] & ~q[1] & ~q[2] & ~q[3]) || 
(~q[0] & q[1] & ~q[2] & ~q[3]) || 
(q[0] & q[1] & ~q[2] & ~q[3]) || 
(~q[0] & ~q[1] & q[2] & ~q[3]) || 
(q[0] & ~q[1] & q[2] & ~q[3]) || 
(~q[0] & q[1] & q[2] & ~q[3]) || 
(q[0] & q[1] & q[2] & ~q[3]) ;

assign r[1] = ~r[0];

assign g[1] = 
(~q[0] & ~q[1] & ~q[2] & ~q[3]) || 
(q[0] & ~q[1] & ~q[2] & ~q[3]) || 
(~q[0] & q[1] & ~q[2] & ~q[3]) || 
(q[0] & q[1] & ~q[2] & ~q[3]) || 
(~q[0] & ~q[1] & q[2] & ~q[3]) || 
(q[0] & ~q[1] & q[2] & ~q[3]) ;
// 8  13
assign g[0] = 
(~q[0] & ~q[1] & ~q[2] & q[3]) || 
(q[0] & ~q[1] & ~q[2] & q[3]) || 
(~q[0] & q[1] & ~q[2] & q[3]) || 
(q[0] & q[1] & ~q[2] & q[3]) || 
(~q[0] & ~q[1] & q[2] & q[3]) || 
(q[0] & ~q[1] & q[2] & q[3]) ;
assign y[1] = 
(~q[0] & q[1] & q[2] & ~q[3]) || 
(q[0] & q[1] & q[2] & ~q[3]) ;
assign y[0] = (~q[0] & q[1] & q[2] & q[3]) || 
(q[0] & q[1] & q[2] & q[3]);


endmodule
